import("EV3_common.cdl");

celltype tTaskMain {
	entry sTaskBody eBody;

};

//[domain(HRP2, "trusted")]
//[domain(HRP2, "nontrusted")]
region rDomainEV3 {
	cell tTaskMain TaskMain {

	};

	cell tTask Task {
	// 呼び口の結合
		cBody = TaskBody.eBody;
		//* 属性の設定
		taskAttribute 	= C_EXP("TA_ACT");
		priority 		= C_EXP("EV3_MRUBY_VM_PRIORITY");
		systemStackSize = C_EXP("MRUBY_VM_STACK_SIZE");
		//userStackSize = C_EXP("STACK_SIZE");
	};

};
