import("EV3_common.cdl");
import("TECSInfo.cdl");
import("tFatFile.cdl");

celltype tTaskMain {
	entry sTaskBody eBody;
	call sLCD cLCD;
	call sButton cButton;
	call sKernel cKernel;
	var {
		int8_t num = 0;
		double64_t num2 = 1.2;
	};
};
// celltype tTemp {
// 	entry sTaskBody eBody;

// 	var {
// 		int8_t dummy = 1;
// 		// int8_t num2;
// 	};
// };
celltype tTECSInfoMain {
	entry sTaskBody	eBody;
	call sLCD cLCD;
	call sButton cButton;
	call sKernel cKernel;
	call sFatFile cFatFile;

  /* TECSInfo */
  call  nTECSInfo::sTECSInfo cTECSInfo;
  [dynamic,optional]
      call  nTECSInfo::sNamespaceInfo cNSInfo;
  [dynamic,optional]
      call  nTECSInfo::sRegionInfo    cRegionInfo;
  [dynamic,optional]
      call  nTECSInfo::sCellInfo      cCellInfo;
  [dynamic,optional]
      call  nTECSInfo::sSignatureInfo cSignatureInfo;
  [dynamic,optional]
      call  nTECSInfo::sCelltypeInfo  cCelltypeInfo;
  [dynamic,optional]
      call  nTECSInfo::sVarDeclInfo   cVarDeclInfo;
  [dynamic,optional]
      call  nTECSInfo::sTypeInfo      cTypeInfo;
  [dynamic,optional]
      call  nTECSInfo::sFunctionInfo  cFunctionInfo;
  [dynamic,optional]
      call  nTECSInfo::sParamInfo     cParamInfo;
  [dynamic,optional]
      call  nTECSInfo::sEntryInfo     cEntryInfo;

  attr {
  	uint8_t BTW = 32;
  	uint8_t NAME_LEN = 32;
  	uint8_t DATA_SIZE = 32;
  };
  var {
  	uint16_t bw;
  	uint16_t num;
  	[size_is(NAME_LEN)]
  		char_t *var_name;
  	[size_is(DATA_SIZE)]
  		char_t *data;
  };
};
//[domain(HRP2, "trusted")]
//[domain(HRP2, "nontrusted")]
region rDomainEV3 {
	// cell tTemp Temp {};

	cell tTaskMain TaskMain {
		cLCD = LCD.eLCD;
		cButton = Button.eButton;
    cKernel = HRP2Kernel.eKernel;
	};
	cell tTask Task {
	// 呼び口の結合
		cBody = TaskMain.eBody;
		// cBody = TECSInfoMain.eBody;
		//* 属性の設定
		taskAttribute 	= C_EXP("TA_ACT");
		priority 		= C_EXP("EV3_MRUBY_VM_PRIORITY");
		systemStackSize = C_EXP("MRUBY_VM_STACK_SIZE");
		//userStackSize = C_EXP("STACK_SIZE");
	};
	/* FatFileセル */
	cell tFatFile FatFile {

	};

	/* TECSInfo */
	cell tTECSInfoMain TECSInfoMain {
    cTECSInfo  = TECSInfo.eTECSInfo;
		cLCD = LCD.eLCD;
		cButton = Button.eButton;
    cKernel = HRP2Kernel.eKernel;
    cFatFile = FatFile.eFatFile;
	};
	cell tCyclicTask TECSInfoTask {
	// 呼び口の結合
		cBody = TECSInfoMain.eBody;
		//* 属性の設定
		cyclicAttribute 	= C_EXP("TA_STA");
		cyclicTime = 100; // 1 = 1msec
		priority = C_EXP("EV3_MRUBY_VM_PRIORITY - 1");
		stackSize = C_EXP("MRUBY_VM_STACK_SIZE"); // systemstacksizeでなくていいのか。kernel.cdlも書き換えなければ
		//userStackSize = C_EXP("STACK_SIZE");
	};
/****** TECSInfo cell ******/
  cell nTECSInfo::tTECSInfo TECSInfo {
      // cTECSInfo = rTECSInfo::TECSInfoSub.eTECSInfo;
      //  この結合は TECSInfoPlugin により生成されるので結合不要
  };
};
